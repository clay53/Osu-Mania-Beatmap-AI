BZh91AY&SY��[ z_�Py����߰?���P>wl�s��ȑB)DmOP�S�i�y�Hz��2 �2Dd)?S�=@  �   	i56���=L�Q�4 �@�A�ɓ&F�L�L))�H�M=Q����2@�@dbd&�r�+b�?ptM*��m�;��� �X���Y [�h� k�+�!vb7�'�(�t(����i�kt�cRBaC�A;霊�F"$LY��Z�@5��ʪ��������d�������iG����t��v�n�����_nǕ��&5�hӫ2���P5���jܪ��8�v������0������2��H:���$��yF�6��cA�"�����Y�η�5i�y�2���w������Vd��r �F�1��*��/�?��M�E�=2�12DD�$�D�P��40�� ��T2��Z�r ��\i9~	Jt��S��'�뜩�����#�f���v�%v�*�e�����ݔ�� ���җtJ�[�#V�r�ddZ�ɽ<����Z[�8�7u�%�Mꊍ�JVH��iû������{�0�Ma�����B�<�f ��,xm��!BU�2D����Z����^k��vF���7�!�M6%jVQ��*)����7_��&�r�o�8����"�!��a�J��8m$w:�jC6vt$'[����x�F�P�@M���H��'+ęb~�]e���F�LGg$<�E6ʠ�0:�M�o, ow��wPnpʻ"��s;�C}�Z	�$<A1�cx$&�75+�#e�8�0:j	X\�؀�B�j�-`(��H�$�	��g;Y[hYhF� y^(��fkY����ř��wC�B� ��٪�n�q�R8�0ߘ3��Ø���C��I����Z��ۆ�6FZ�a8�&5kCN�v\�4�T����<�6���@^���[��bᠬveX����,��

Ʒ�L�{JK)t�tk���x��R��51��!ndk���"�(Hx~-�